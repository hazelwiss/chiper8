`timescale 1ns/100ps

`define TRUE 1'b1
`define FALSE 1'b0