`include "verilog/include/defs.sv"

module dcache();

endmodule 